
module dec_test (
	clk_clk,
	reset_reset_n,
	sem_export_train,
	sem_export_red,
	sem_export_yellow,
	sem_export_green);	

	input		clk_clk;
	input		reset_reset_n;
	input		sem_export_train;
	output		sem_export_red;
	output		sem_export_yellow;
	output		sem_export_green;
endmodule
