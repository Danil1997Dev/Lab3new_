`timescale 1ps / 1ps

module tb ();

   dec_test_tb dut();
   test_program tp();

endmodule 
