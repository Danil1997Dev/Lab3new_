// dec_test_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module dec_test_tb (
	);

	wire        dec_test_inst_clk_bfm_clk_clk;              // dec_test_inst_clk_bfm:clk -> [dec_test_inst:clk_clk, dec_test_inst_reset_bfm:clk]
	wire        dec_test_inst_sem_export_red;               // dec_test_inst:sem_export_red -> dec_test_inst_sem_export_bfm:sig_red
	wire        dec_test_inst_sem_export_green;             // dec_test_inst:sem_export_green -> dec_test_inst_sem_export_bfm:sig_green
	wire        dec_test_inst_sem_export_yellow;            // dec_test_inst:sem_export_yellow -> dec_test_inst_sem_export_bfm:sig_yellow
	wire  [0:0] dec_test_inst_sem_export_bfm_conduit_train; // dec_test_inst_sem_export_bfm:sig_train -> dec_test_inst:sem_export_train
	wire        dec_test_inst_reset_bfm_reset_reset;        // dec_test_inst_reset_bfm:reset -> dec_test_inst:reset_reset_n

	dec_test dec_test_inst (
		.clk_clk           (dec_test_inst_clk_bfm_clk_clk),              //        clk.clk
		.reset_reset_n     (dec_test_inst_reset_bfm_reset_reset),        //      reset.reset_n
		.sem_export_train  (dec_test_inst_sem_export_bfm_conduit_train), // sem_export.train
		.sem_export_red    (dec_test_inst_sem_export_red),               //           .red
		.sem_export_yellow (dec_test_inst_sem_export_yellow),            //           .yellow
		.sem_export_green  (dec_test_inst_sem_export_green)              //           .green
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) dec_test_inst_clk_bfm (
		.clk (dec_test_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) dec_test_inst_reset_bfm (
		.reset (dec_test_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (dec_test_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm dec_test_inst_sem_export_bfm (
		.sig_green  (dec_test_inst_sem_export_green),             // conduit.green
		.sig_red    (dec_test_inst_sem_export_red),               //        .red
		.sig_train  (dec_test_inst_sem_export_bfm_conduit_train), //        .train
		.sig_yellow (dec_test_inst_sem_export_yellow)             //        .yellow
	);

endmodule
